magic
tech sky130A
magscale 1 2
timestamp 1745519855
<< checkpaint >>
rect -3932 -2564 9766 13580
<< viali >>
rect 2237 9129 2271 9163
rect 1869 9061 1903 9095
rect 1685 8925 1719 8959
rect 2053 8925 2087 8959
rect 2421 8925 2455 8959
rect 1501 8789 1535 8823
rect 1685 8449 1719 8483
rect 4077 8449 4111 8483
rect 4537 8449 4571 8483
rect 4215 8381 4249 8415
rect 1501 8313 1535 8347
rect 4353 8245 4387 8279
rect 4445 8245 4479 8279
rect 2329 7905 2363 7939
rect 2789 7905 2823 7939
rect 4353 7905 4387 7939
rect 1685 7837 1719 7871
rect 2697 7837 2731 7871
rect 4537 7837 4571 7871
rect 5181 7837 5215 7871
rect 5365 7837 5399 7871
rect 5273 7769 5307 7803
rect 1501 7701 1535 7735
rect 4721 7701 4755 7735
rect 3249 7497 3283 7531
rect 1685 7361 1719 7395
rect 3157 7361 3191 7395
rect 3341 7361 3375 7395
rect 5457 7361 5491 7395
rect 1501 7157 1535 7191
rect 5273 7157 5307 7191
rect 1685 6749 1719 6783
rect 1501 6613 1535 6647
rect 1685 6273 1719 6307
rect 1869 6273 1903 6307
rect 2145 6273 2179 6307
rect 1961 6137 1995 6171
rect 2053 6137 2087 6171
rect 1501 6069 1535 6103
rect 2329 6069 2363 6103
rect 1409 5661 1443 5695
rect 1593 5525 1627 5559
rect 2789 5253 2823 5287
rect 1409 5185 1443 5219
rect 3065 5185 3099 5219
rect 2881 5117 2915 5151
rect 1593 5049 1627 5083
rect 2421 5049 2455 5083
rect 2329 4981 2363 5015
rect 3249 4981 3283 5015
rect 3433 4777 3467 4811
rect 4445 4777 4479 4811
rect 4905 4777 4939 4811
rect 2697 4709 2731 4743
rect 3801 4709 3835 4743
rect 2973 4641 3007 4675
rect 4261 4641 4295 4675
rect 1409 4573 1443 4607
rect 3065 4573 3099 4607
rect 3433 4573 3467 4607
rect 3617 4573 3651 4607
rect 4169 4573 4203 4607
rect 4629 4573 4663 4607
rect 4721 4573 4755 4607
rect 4445 4505 4479 4539
rect 1593 4437 1627 4471
rect 1593 4233 1627 4267
rect 1409 4097 1443 4131
rect 2421 4097 2455 4131
rect 2605 4097 2639 4131
rect 2605 3961 2639 3995
rect 1777 3689 1811 3723
rect 1409 3485 1443 3519
rect 1961 3485 1995 3519
rect 1593 3349 1627 3383
rect 3433 3145 3467 3179
rect 5457 3145 5491 3179
rect 4997 3077 5031 3111
rect 1777 3009 1811 3043
rect 3617 3009 3651 3043
rect 5273 3009 5307 3043
rect 1593 2941 1627 2975
rect 5089 2941 5123 2975
rect 1961 2873 1995 2907
rect 4997 2805 5031 2839
rect 2145 2601 2179 2635
rect 1869 2533 1903 2567
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 1961 2397 1995 2431
rect 1593 2261 1627 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 1302 9120 1308 9172
rect 1360 9160 1366 9172
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 1360 9132 2237 9160
rect 1360 9120 1366 9132
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 2225 9123 2283 9129
rect 934 9052 940 9104
rect 992 9092 998 9104
rect 1857 9095 1915 9101
rect 1857 9092 1869 9095
rect 992 9064 1869 9092
rect 992 9052 998 9064
rect 1857 9061 1869 9064
rect 1903 9061 1915 9095
rect 1857 9055 1915 9061
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 1854 8956 1860 8968
rect 1719 8928 1860 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2409 8959 2467 8965
rect 2409 8925 2421 8959
rect 2455 8956 2467 8959
rect 3326 8956 3332 8968
rect 2455 8928 3332 8956
rect 2455 8925 2467 8928
rect 2409 8919 2467 8925
rect 2056 8888 2084 8919
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 3050 8888 3056 8900
rect 2056 8860 3056 8888
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 842 8780 848 8832
rect 900 8820 906 8832
rect 1489 8823 1547 8829
rect 1489 8820 1501 8823
rect 900 8792 1501 8820
rect 900 8780 906 8792
rect 1489 8789 1501 8792
rect 1535 8789 1547 8823
rect 1489 8783 1547 8789
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3200 8452 4077 8480
rect 3200 8440 3206 8452
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 5074 8480 5080 8492
rect 4571 8452 5080 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 4203 8415 4261 8421
rect 4203 8381 4215 8415
rect 4249 8412 4261 8415
rect 4338 8412 4344 8424
rect 4249 8384 4344 8412
rect 4249 8381 4261 8384
rect 4203 8375 4261 8381
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4341 8279 4399 8285
rect 4341 8276 4353 8279
rect 4212 8248 4353 8276
rect 4212 8236 4218 8248
rect 4341 8245 4353 8248
rect 4387 8245 4399 8279
rect 4341 8239 4399 8245
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4522 8276 4528 8288
rect 4479 8248 4528 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 1762 7896 1768 7948
rect 1820 7936 1826 7948
rect 2317 7939 2375 7945
rect 2317 7936 2329 7939
rect 1820 7908 2329 7936
rect 1820 7896 1826 7908
rect 2317 7905 2329 7908
rect 2363 7905 2375 7939
rect 2317 7899 2375 7905
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 2823 7908 4353 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 4341 7905 4353 7908
rect 4387 7936 4399 7939
rect 4430 7936 4436 7948
rect 4387 7908 4436 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1688 7800 1716 7831
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 2685 7871 2743 7877
rect 2685 7868 2697 7871
rect 2464 7840 2697 7868
rect 2464 7828 2470 7840
rect 2685 7837 2697 7840
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 1688 7772 5273 7800
rect 5261 7769 5273 7772
rect 5307 7769 5319 7803
rect 5261 7763 5319 7769
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 1489 7735 1547 7741
rect 1489 7732 1501 7735
rect 900 7704 1501 7732
rect 900 7692 906 7704
rect 1489 7701 1501 7704
rect 1535 7701 1547 7735
rect 1489 7695 1547 7701
rect 4706 7692 4712 7744
rect 4764 7692 4770 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 3237 7531 3295 7537
rect 3237 7497 3249 7531
rect 3283 7528 3295 7531
rect 4246 7528 4252 7540
rect 3283 7500 4252 7528
rect 3283 7497 3295 7500
rect 3237 7491 3295 7497
rect 4246 7488 4252 7500
rect 4304 7528 4310 7540
rect 5350 7528 5356 7540
rect 4304 7500 5356 7528
rect 4304 7488 4310 7500
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1688 7324 1716 7355
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7392 3387 7395
rect 4154 7392 4160 7404
rect 3375 7364 4160 7392
rect 3375 7361 3387 7364
rect 3329 7355 3387 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4706 7352 4712 7404
rect 4764 7392 4770 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 4764 7364 5457 7392
rect 4764 7352 4770 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 3786 7324 3792 7336
rect 1688 7296 3792 7324
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 5258 7148 5264 7200
rect 5316 7148 5322 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 5258 6780 5264 6792
rect 1719 6752 5264 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 1210 6604 1216 6656
rect 1268 6644 1274 6656
rect 1489 6647 1547 6653
rect 1489 6644 1501 6647
rect 1268 6616 1501 6644
rect 1268 6604 1274 6616
rect 1489 6613 1501 6616
rect 1535 6613 1547 6647
rect 1489 6607 1547 6613
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 1762 6304 1768 6316
rect 1719 6276 1768 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6304 2191 6307
rect 2498 6304 2504 6316
rect 2179 6276 2504 6304
rect 2179 6273 2191 6276
rect 2133 6267 2191 6273
rect 1578 6196 1584 6248
rect 1636 6236 1642 6248
rect 1872 6236 1900 6267
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 1636 6208 1900 6236
rect 1636 6196 1642 6208
rect 1762 6128 1768 6180
rect 1820 6168 1826 6180
rect 1949 6171 2007 6177
rect 1949 6168 1961 6171
rect 1820 6140 1961 6168
rect 1820 6128 1826 6140
rect 1949 6137 1961 6140
rect 1995 6137 2007 6171
rect 1949 6131 2007 6137
rect 2041 6171 2099 6177
rect 2041 6137 2053 6171
rect 2087 6168 2099 6171
rect 3142 6168 3148 6180
rect 2087 6140 3148 6168
rect 2087 6137 2099 6140
rect 2041 6131 2099 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 842 6060 848 6112
rect 900 6100 906 6112
rect 1489 6103 1547 6109
rect 1489 6100 1501 6103
rect 900 6072 1501 6100
rect 900 6060 906 6072
rect 1489 6069 1501 6072
rect 1535 6069 1547 6103
rect 1489 6063 1547 6069
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2958 6100 2964 6112
rect 2363 6072 2964 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 3142 5556 3148 5568
rect 1627 5528 3148 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 2777 5287 2835 5293
rect 2777 5253 2789 5287
rect 2823 5284 2835 5287
rect 2958 5284 2964 5296
rect 2823 5256 2964 5284
rect 2823 5253 2835 5256
rect 2777 5247 2835 5253
rect 2958 5244 2964 5256
rect 3016 5244 3022 5296
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 3142 5216 3148 5228
rect 3099 5188 3148 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 2498 5148 2504 5160
rect 1596 5120 2504 5148
rect 1596 5089 1624 5120
rect 2498 5108 2504 5120
rect 2556 5148 2562 5160
rect 2869 5151 2927 5157
rect 2869 5148 2881 5151
rect 2556 5120 2881 5148
rect 2556 5108 2562 5120
rect 2869 5117 2881 5120
rect 2915 5148 2927 5151
rect 4706 5148 4712 5160
rect 2915 5120 4712 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5049 1639 5083
rect 2409 5083 2467 5089
rect 2409 5080 2421 5083
rect 1581 5043 1639 5049
rect 2240 5052 2421 5080
rect 1486 4972 1492 5024
rect 1544 5012 1550 5024
rect 2240 5012 2268 5052
rect 2409 5049 2421 5052
rect 2455 5080 2467 5083
rect 4154 5080 4160 5092
rect 2455 5052 4160 5080
rect 2455 5049 2467 5052
rect 2409 5043 2467 5049
rect 4154 5040 4160 5052
rect 4212 5080 4218 5092
rect 4890 5080 4896 5092
rect 4212 5052 4896 5080
rect 4212 5040 4218 5052
rect 4890 5040 4896 5052
rect 4948 5040 4954 5092
rect 1544 4984 2268 5012
rect 1544 4972 1550 4984
rect 2314 4972 2320 5024
rect 2372 4972 2378 5024
rect 3237 5015 3295 5021
rect 3237 4981 3249 5015
rect 3283 5012 3295 5015
rect 3418 5012 3424 5024
rect 3283 4984 3424 5012
rect 3283 4981 3295 4984
rect 3237 4975 3295 4981
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 3050 4768 3056 4820
rect 3108 4808 3114 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 3108 4780 3433 4808
rect 3108 4768 3114 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 3421 4771 3479 4777
rect 3528 4780 4445 4808
rect 1854 4700 1860 4752
rect 1912 4740 1918 4752
rect 2685 4743 2743 4749
rect 2685 4740 2697 4743
rect 1912 4712 2697 4740
rect 1912 4700 1918 4712
rect 2685 4709 2697 4712
rect 2731 4709 2743 4743
rect 2685 4703 2743 4709
rect 3142 4700 3148 4752
rect 3200 4740 3206 4752
rect 3528 4740 3556 4780
rect 4433 4777 4445 4780
rect 4479 4777 4491 4811
rect 4433 4771 4491 4777
rect 4890 4768 4896 4820
rect 4948 4768 4954 4820
rect 3200 4712 3556 4740
rect 3200 4700 3206 4712
rect 3786 4700 3792 4752
rect 3844 4700 3850 4752
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 3016 4644 3648 4672
rect 3016 4632 3022 4644
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 1762 4536 1768 4548
rect 1596 4508 1768 4536
rect 1596 4477 1624 4508
rect 1762 4496 1768 4508
rect 1820 4536 1826 4548
rect 3068 4536 3096 4567
rect 3418 4564 3424 4616
rect 3476 4564 3482 4616
rect 3620 4613 3648 4644
rect 4246 4632 4252 4684
rect 4304 4632 4310 4684
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 4264 4576 4629 4604
rect 4264 4536 4292 4576
rect 4617 4573 4629 4576
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 1820 4508 4292 4536
rect 4433 4539 4491 4545
rect 1820 4496 1826 4508
rect 4433 4505 4445 4539
rect 4479 4505 4491 4539
rect 4433 4499 4491 4505
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4437 1639 4471
rect 1581 4431 1639 4437
rect 1854 4428 1860 4480
rect 1912 4468 1918 4480
rect 4448 4468 4476 4499
rect 1912 4440 4476 4468
rect 1912 4428 1918 4440
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 1578 4224 1584 4276
rect 1636 4264 1642 4276
rect 1854 4264 1860 4276
rect 1636 4236 1860 4264
rect 1636 4224 1642 4236
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 992 4100 1409 4128
rect 992 4088 998 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2498 4128 2504 4140
rect 2455 4100 2504 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 3142 4128 3148 4140
rect 2639 4100 3148 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 3142 4088 3148 4100
rect 3200 4128 3206 4140
rect 3602 4128 3608 4140
rect 3200 4100 3608 4128
rect 3200 4088 3206 4100
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 2593 3995 2651 4001
rect 2593 3961 2605 3995
rect 2639 3992 2651 3995
rect 2958 3992 2964 4004
rect 2639 3964 2964 3992
rect 2639 3961 2651 3964
rect 2593 3955 2651 3961
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 1765 3723 1823 3729
rect 1765 3720 1777 3723
rect 1728 3692 1777 3720
rect 1728 3680 1734 3692
rect 1765 3689 1777 3692
rect 1811 3689 1823 3723
rect 1765 3683 1823 3689
rect 842 3476 848 3528
rect 900 3516 906 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 900 3488 1409 3516
rect 900 3476 906 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3516 2007 3519
rect 2314 3516 2320 3528
rect 1995 3488 2320 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 1578 3340 1584 3392
rect 1636 3340 1642 3392
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3421 3179 3479 3185
rect 3421 3176 3433 3179
rect 3384 3148 3433 3176
rect 3384 3136 3390 3148
rect 3421 3145 3433 3148
rect 3467 3145 3479 3179
rect 3421 3139 3479 3145
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 4488 3148 5457 3176
rect 4488 3136 4494 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5445 3139 5503 3145
rect 4890 3068 4896 3120
rect 4948 3108 4954 3120
rect 4985 3111 5043 3117
rect 4985 3108 4997 3111
rect 4948 3080 4997 3108
rect 4948 3068 4954 3080
rect 4985 3077 4997 3080
rect 5031 3077 5043 3111
rect 4985 3071 5043 3077
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1544 3012 1777 3040
rect 1544 3000 1550 3012
rect 1765 3009 1777 3012
rect 1811 3009 1823 3043
rect 1765 3003 1823 3009
rect 3602 3000 3608 3052
rect 3660 3000 3666 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 3712 3012 5273 3040
rect 1578 2932 1584 2984
rect 1636 2972 1642 2984
rect 3234 2972 3240 2984
rect 1636 2944 3240 2972
rect 1636 2932 1642 2944
rect 3234 2932 3240 2944
rect 3292 2972 3298 2984
rect 3712 2972 3740 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 3292 2944 3740 2972
rect 3292 2932 3298 2944
rect 5074 2932 5080 2984
rect 5132 2932 5138 2984
rect 1949 2907 2007 2913
rect 1949 2873 1961 2907
rect 1995 2904 2007 2907
rect 5166 2904 5172 2916
rect 1995 2876 5172 2904
rect 1995 2873 2007 2876
rect 1949 2867 2007 2873
rect 5166 2864 5172 2876
rect 5224 2864 5230 2916
rect 4982 2796 4988 2848
rect 5040 2796 5046 2848
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 2406 2632 2412 2644
rect 2179 2604 2412 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 1857 2567 1915 2573
rect 1857 2533 1869 2567
rect 1903 2564 1915 2567
rect 5074 2564 5080 2576
rect 1903 2536 5080 2564
rect 1903 2533 1915 2536
rect 1857 2527 1915 2533
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 1026 2456 1032 2508
rect 1084 2496 1090 2508
rect 1084 2468 1992 2496
rect 1084 2456 1090 2468
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1964 2437 1992 2468
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 934 2320 940 2372
rect 992 2360 998 2372
rect 1688 2360 1716 2391
rect 992 2332 1716 2360
rect 992 2320 998 2332
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 4154 2292 4160 2304
rect 1627 2264 4160 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 4154 2252 4160 2264
rect 4212 2292 4218 2304
rect 4982 2292 4988 2304
rect 4212 2264 4988 2292
rect 4212 2252 4218 2264
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 1308 9120 1360 9172
rect 940 9052 992 9104
rect 1860 8916 1912 8968
rect 3332 8916 3384 8968
rect 3056 8848 3108 8900
rect 848 8780 900 8832
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 3148 8440 3200 8492
rect 5080 8440 5132 8492
rect 4344 8372 4396 8424
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 4160 8236 4212 8288
rect 4528 8236 4580 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 1768 7896 1820 7948
rect 4436 7896 4488 7948
rect 2412 7828 2464 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 848 7692 900 7744
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 4252 7488 4304 7540
rect 5356 7488 5408 7540
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 4160 7352 4212 7404
rect 4712 7352 4764 7404
rect 3792 7284 3844 7336
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 5264 6740 5316 6792
rect 1216 6604 1268 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 1768 6264 1820 6316
rect 1584 6196 1636 6248
rect 2504 6264 2556 6316
rect 1768 6128 1820 6180
rect 3148 6128 3200 6180
rect 848 6060 900 6112
rect 2964 6060 3016 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 3148 5516 3200 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 2964 5244 3016 5296
rect 848 5176 900 5228
rect 3148 5176 3200 5228
rect 2504 5108 2556 5160
rect 4712 5108 4764 5160
rect 1492 4972 1544 5024
rect 4160 5040 4212 5092
rect 4896 5040 4948 5092
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 3424 4972 3476 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 3056 4768 3108 4820
rect 1860 4700 1912 4752
rect 3148 4700 3200 4752
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 3792 4743 3844 4752
rect 3792 4709 3801 4743
rect 3801 4709 3835 4743
rect 3835 4709 3844 4743
rect 3792 4700 3844 4709
rect 2964 4675 3016 4684
rect 2964 4641 2973 4675
rect 2973 4641 3007 4675
rect 3007 4641 3016 4675
rect 2964 4632 3016 4641
rect 848 4564 900 4616
rect 1768 4496 1820 4548
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 1860 4428 1912 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 1860 4224 1912 4276
rect 940 4088 992 4140
rect 2504 4088 2556 4140
rect 3148 4088 3200 4140
rect 3608 4088 3660 4140
rect 2964 3952 3016 4004
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 1676 3680 1728 3732
rect 848 3476 900 3528
rect 2320 3476 2372 3528
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 3332 3136 3384 3188
rect 4436 3136 4488 3188
rect 4896 3068 4948 3120
rect 1492 3000 1544 3052
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 3240 2932 3292 2984
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 5172 2864 5224 2916
rect 4988 2839 5040 2848
rect 4988 2805 4997 2839
rect 4997 2805 5031 2839
rect 5031 2805 5040 2839
rect 4988 2796 5040 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 2412 2592 2464 2644
rect 5080 2524 5132 2576
rect 1032 2456 1084 2508
rect 848 2388 900 2440
rect 940 2320 992 2372
rect 4160 2252 4212 2304
rect 4988 2252 5040 2304
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1306 9616 1362 9625
rect 1306 9551 1362 9560
rect 1320 9178 1348 9551
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 940 9104 992 9110
rect 938 9072 940 9081
rect 992 9072 994 9081
rect 938 9007 994 9016
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 848 8832 900 8838
rect 848 8774 900 8780
rect 860 8673 888 8774
rect 846 8664 902 8673
rect 846 8599 902 8608
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 7993 1532 8298
rect 1490 7984 1546 7993
rect 1490 7919 1546 7928
rect 848 7744 900 7750
rect 848 7686 900 7692
rect 860 7585 888 7686
rect 846 7576 902 7585
rect 846 7511 902 7520
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1216 6656 1268 6662
rect 1216 6598 1268 6604
rect 1228 6361 1256 6598
rect 1214 6352 1270 6361
rect 1214 6287 1270 6296
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 848 6112 900 6118
rect 848 6054 900 6060
rect 860 5953 888 6054
rect 846 5944 902 5953
rect 846 5879 902 5888
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5273 1440 5646
rect 1398 5264 1454 5273
rect 848 5228 900 5234
rect 1398 5199 1454 5208
rect 848 5170 900 5176
rect 860 4865 888 5170
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 846 4856 902 4865
rect 846 4791 902 4800
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 860 4321 888 4558
rect 846 4312 902 4321
rect 846 4247 902 4256
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 3641 980 4082
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 848 3528 900 3534
rect 848 3470 900 3476
rect 860 3233 888 3470
rect 846 3224 902 3233
rect 846 3159 902 3168
rect 1504 3058 1532 4966
rect 1596 4282 1624 6190
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1688 3738 1716 8434
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1780 6322 1808 7890
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1780 4554 1808 6122
rect 1872 4758 1900 8910
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1860 4752 1912 4758
rect 1860 4694 1912 4700
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4282 1900 4422
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 2332 3534 2360 4966
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1596 2990 1624 3334
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2424 2650 2452 7822
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2516 5166 2544 6258
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2976 5302 3004 6054
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2516 4146 2544 5102
rect 3068 4826 3096 8842
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3160 7410 3188 8434
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 6914 3188 7346
rect 3160 6886 3280 6914
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3160 5574 3188 6122
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3160 5234 3188 5510
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3160 4758 3188 5170
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2976 4010 3004 4626
rect 3160 4146 3188 4694
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 3252 2990 3280 6886
rect 3344 3194 3372 8910
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 7410 4200 8230
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3436 4622 3464 4966
rect 3804 4758 3832 7278
rect 4172 5098 4200 7346
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 4264 4690 4292 7482
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 4160 4616 4212 4622
rect 4356 4570 4384 8366
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4212 4564 4384 4570
rect 4160 4558 4384 4564
rect 4172 4542 4384 4558
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3620 3058 3648 4082
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 1032 2508 1084 2514
rect 1032 2450 1084 2456
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 900 2408 902 2417
rect 846 2343 902 2352
rect 940 2372 992 2378
rect 940 2314 992 2320
rect 952 2009 980 2314
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 1044 1465 1072 2450
rect 4172 2310 4200 4542
rect 4448 3194 4476 7890
rect 4540 7886 4568 8230
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4724 7410 4752 7686
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4724 4622 4752 5102
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4908 4826 4936 5034
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4908 3126 4936 4762
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 5092 2990 5120 8434
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 5000 2310 5028 2790
rect 5092 2582 5120 2926
rect 5184 2922 5212 7822
rect 5368 7546 5396 7822
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6798 5304 7142
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 1030 1456 1086 1465
rect 1030 1391 1086 1400
<< via2 >>
rect 1306 9560 1362 9616
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 938 9052 940 9072
rect 940 9052 992 9072
rect 992 9052 994 9072
rect 938 9016 994 9052
rect 846 8608 902 8664
rect 1490 7928 1546 7984
rect 846 7520 902 7576
rect 1490 6840 1546 6896
rect 1214 6296 1270 6352
rect 846 5888 902 5944
rect 1398 5208 1454 5264
rect 846 4800 902 4856
rect 846 4256 902 4312
rect 938 3576 994 3632
rect 846 3168 902 3224
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 938 1944 994 2000
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1030 1400 1086 1456
<< metal3 >>
rect 0 9618 800 9648
rect 1301 9618 1367 9621
rect 0 9616 1367 9618
rect 0 9560 1306 9616
rect 1362 9560 1367 9616
rect 0 9558 1367 9560
rect 0 9528 800 9558
rect 1301 9555 1367 9558
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 841 8666 907 8669
rect 798 8664 907 8666
rect 798 8608 846 8664
rect 902 8608 907 8664
rect 798 8603 907 8608
rect 798 8560 858 8603
rect 0 8470 858 8560
rect 0 8440 800 8470
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 0 7986 800 8016
rect 1485 7986 1551 7989
rect 0 7984 1551 7986
rect 0 7928 1490 7984
rect 1546 7928 1551 7984
rect 0 7926 1551 7928
rect 0 7896 800 7926
rect 1485 7923 1551 7926
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 841 7578 907 7581
rect 798 7576 907 7578
rect 798 7520 846 7576
rect 902 7520 907 7576
rect 798 7515 907 7520
rect 798 7472 858 7515
rect 0 7382 858 7472
rect 0 7352 800 7382
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 0 6354 800 6384
rect 1209 6354 1275 6357
rect 0 6352 1275 6354
rect 0 6296 1214 6352
rect 1270 6296 1275 6352
rect 0 6294 1275 6296
rect 0 6264 800 6294
rect 1209 6291 1275 6294
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 841 5946 907 5949
rect 798 5944 907 5946
rect 798 5888 846 5944
rect 902 5888 907 5944
rect 798 5883 907 5888
rect 798 5840 858 5883
rect 0 5750 858 5840
rect 0 5720 800 5750
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 0 5266 800 5296
rect 1393 5266 1459 5269
rect 0 5264 1459 5266
rect 0 5208 1398 5264
rect 1454 5208 1459 5264
rect 0 5206 1459 5208
rect 0 5176 800 5206
rect 1393 5203 1459 5206
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 841 4858 907 4861
rect 798 4856 907 4858
rect 798 4800 846 4856
rect 902 4800 907 4856
rect 798 4795 907 4800
rect 798 4752 858 4795
rect 0 4662 858 4752
rect 0 4632 800 4662
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 841 4314 907 4317
rect 798 4312 907 4314
rect 798 4256 846 4312
rect 902 4256 907 4312
rect 798 4251 907 4256
rect 798 4208 858 4251
rect 0 4118 858 4208
rect 0 4088 800 4118
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 841 3226 907 3229
rect 798 3224 907 3226
rect 798 3168 846 3224
rect 902 3168 907 3224
rect 798 3163 907 3168
rect 798 3120 858 3163
rect 0 3030 858 3120
rect 0 3000 800 3030
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 0 2546 800 2576
rect 0 2456 858 2546
rect 798 2413 858 2456
rect 798 2408 907 2413
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2350 907 2352
rect 841 2347 907 2350
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
rect 0 1458 800 1488
rect 1025 1458 1091 1461
rect 0 1456 1091 1458
rect 0 1400 1030 1456
rect 1086 1400 1091 1456
rect 0 1398 1091 1400
rect 0 1368 800 1398
rect 1025 1395 1091 1398
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform -1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _11_
timestamp 0
transform -1 0 3312 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _12_
timestamp 0
transform -1 0 2392 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _13_
timestamp 0
transform 1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _14_
timestamp 0
transform -1 0 2852 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 0
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _16_
timestamp 0
transform -1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _17_
timestamp 0
transform 1 0 1564 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _19_
timestamp 0
transform -1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _20_
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _21_
timestamp 0
transform 1 0 4048 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform 1 0 4324 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _24_
timestamp 0
transform -1 0 2944 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _25_
timestamp 0
transform 1 0 2852 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _26_
timestamp 0
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 0
transform 1 0 3404 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_12
timestamp 0
transform 1 0 2208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_24
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_47
timestamp 0
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_10
timestamp 0
transform 1 0 2024 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_22
timestamp 0
transform 1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_28
timestamp 0
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_40
timestamp 0
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_6
timestamp 0
transform 1 0 1656 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_10
timestamp 0
transform 1 0 2024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_22
timestamp 0
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 0
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_6
timestamp 0
transform 1 0 1656 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_17
timestamp 0
transform 1 0 2668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_29
timestamp 0
transform 1 0 3772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_41
timestamp 0
transform 1 0 4876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_47
timestamp 0
transform 1 0 5428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_6
timestamp 0
transform 1 0 1656 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_14
timestamp 0
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_24
timestamp 0
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_43
timestamp 0
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_6
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_12
timestamp 0
transform 1 0 2208 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_24
timestamp 0
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_36
timestamp 0
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 0
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_14
timestamp 0
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_26
timestamp 0
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_38
timestamp 0
transform 1 0 4600 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_46
timestamp 0
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_7
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_19
timestamp 0
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_47
timestamp 0
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_7
timestamp 0
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_19
timestamp 0
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_25
timestamp 0
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_37
timestamp 0
transform 1 0 4508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_7
timestamp 0
transform 1 0 1748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_20
timestamp 0
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_40
timestamp 0
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_47
timestamp 0
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_7
timestamp 0
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_19
timestamp 0
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_31
timestamp 0
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_38
timestamp 0
transform 1 0 4600 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_46
timestamp 0
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_47
timestamp 0
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform -1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform -1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
rlabel metal1 s 3450 8704 3450 8704 4 VGND
rlabel metal1 s 3450 9248 3450 9248 4 VPWR
rlabel metal2 s 2990 4318 2990 4318 4 _00_
rlabel metal1 s 2898 5270 2898 5270 4 _01_
rlabel metal1 s 2346 5066 2346 5066 4 _02_
rlabel metal1 s 2162 3502 2162 3502 4 _03_
rlabel metal1 s 4324 7514 4324 7514 4 _04_
rlabel metal1 s 3588 2890 3588 2890 4 _05_
rlabel metal1 s 4968 3162 4968 3162 4 _06_
rlabel metal2 s 4554 8058 4554 8058 4 _07_
rlabel metal1 s 5106 7378 5106 7378 4 _08_
rlabel metal2 s 3450 4794 3450 4794 4 _09_
rlabel metal3 s 1050 5236 1050 5236 4 a1[0]
rlabel metal3 s 0 4632 800 4752 4 a1[1]
port 4 nsew
rlabel metal3 s 0 4088 800 4208 4 a1[2]
port 5 nsew
rlabel metal3 s 820 3604 820 3604 4 a1[3]
rlabel metal3 s 0 3000 800 3120 4 a1[4]
port 7 nsew
rlabel metal3 s 0 2456 800 2576 4 a1[5]
port 8 nsew
rlabel metal3 s 820 1972 820 1972 4 a1[6]
rlabel metal3 s 866 1428 866 1428 4 a1[7]
rlabel metal1 s 1794 9146 1794 9146 4 b1[0]
rlabel metal3 s 820 9044 820 9044 4 b1[1]
rlabel metal3 s 0 8440 800 8560 4 b1[2]
port 13 nsew
rlabel metal3 s 1096 7956 1096 7956 4 b1[3]
rlabel metal3 s 0 7352 800 7472 4 b1[4]
port 15 nsew
rlabel metal3 s 1096 6868 1096 6868 4 b1[5]
rlabel metal1 s 1380 6630 1380 6630 4 b1[6]
rlabel metal3 s 0 5720 800 5840 4 b1[7]
port 18 nsew
rlabel metal1 s 3128 4114 3128 4114 4 net1
rlabel metal1 s 3266 4794 3266 4794 4 net10
rlabel metal1 s 2300 4726 2300 4726 4 net11
rlabel metal1 s 1748 3706 1748 3706 4 net12
rlabel metal1 s 1702 7820 1702 7820 4 net13
rlabel metal1 s 2760 7310 2760 7310 4 net14
rlabel metal1 s 3496 6766 3496 6766 4 net15
rlabel metal1 s 1748 6290 1748 6290 4 net16
rlabel metal1 s 3818 5134 3818 5134 4 net2
rlabel metal1 s 3082 4556 3082 4556 4 net3
rlabel metal1 s 1748 4250 1748 4250 4 net4
rlabel metal1 s 2668 2958 2668 2958 4 net5
rlabel metal2 s 5014 2550 5014 2550 4 net6
rlabel metal1 s 3496 2550 3496 2550 4 net7
rlabel metal1 s 2300 2618 2300 2618 4 net8
rlabel metal1 s 3404 3162 3404 3162 4 net9
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 5176 800 5296 0 FreeSans 600 0 0 0 a1[0]
port 3 nsew
flabel metal3 s 400 4692 400 4692 0 FreeSans 600 0 0 0 a1[1]
flabel metal3 s 400 4148 400 4148 0 FreeSans 600 0 0 0 a1[2]
flabel metal3 s 0 3544 800 3664 0 FreeSans 600 0 0 0 a1[3]
port 6 nsew
flabel metal3 s 400 3060 400 3060 0 FreeSans 600 0 0 0 a1[4]
flabel metal3 s 400 2516 400 2516 0 FreeSans 600 0 0 0 a1[5]
flabel metal3 s 0 1912 800 2032 0 FreeSans 600 0 0 0 a1[6]
port 9 nsew
flabel metal3 s 0 1368 800 1488 0 FreeSans 600 0 0 0 a1[7]
port 10 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 b1[0]
port 11 nsew
flabel metal3 s 0 8984 800 9104 0 FreeSans 600 0 0 0 b1[1]
port 12 nsew
flabel metal3 s 400 8500 400 8500 0 FreeSans 600 0 0 0 b1[2]
flabel metal3 s 0 7896 800 8016 0 FreeSans 600 0 0 0 b1[3]
port 14 nsew
flabel metal3 s 400 7412 400 7412 0 FreeSans 600 0 0 0 b1[4]
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 b1[5]
port 16 nsew
flabel metal3 s 0 6264 800 6384 0 FreeSans 600 0 0 0 b1[6]
port 17 nsew
flabel metal3 s 400 5780 400 5780 0 FreeSans 600 0 0 0 b1[7]
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
