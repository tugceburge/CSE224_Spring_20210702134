* NGSPICE file created from twos_complement.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt twos_complement VGND VPWR a1[0] a1[1] a1[2] a1[3] a1[4] a1[5] a1[6] a1[7]
+ b1[0] b1[1] b1[2] b1[3] b1[4] b1[5] b1[6] b1[7]
XTAP_TAPCELL_ROW_12_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput10 net10 VGND VGND VPWR VPWR b1[1] sky130_fd_sc_hd__buf_2
XFILLER_0_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput9 net9 VGND VGND VPWR VPWR b1[0] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR b1[2] sky130_fd_sc_hd__buf_2
XFILLER_0_11_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput12 net12 VGND VGND VPWR VPWR b1[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput13 net13 VGND VGND VPWR VPWR b1[4] sky130_fd_sc_hd__buf_2
XFILLER_0_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27_ net1 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
Xoutput14 net14 VGND VGND VPWR VPWR b1[5] sky130_fd_sc_hd__buf_2
XFILLER_0_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26_ _00_ _09_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR b1[6] sky130_fd_sc_hd__buf_2
XFILLER_0_9_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25_ net2 net1 VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__and2_1
Xoutput16 net16 VGND VGND VPWR VPWR b1[7] sky130_fd_sc_hd__buf_2
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24_ net8 _06_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_11_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23_ _08_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22_ _06_ _07_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21_ net5 net6 _02_ net7 VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_1_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20_ net5 net6 net7 _02_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__or4_1
Xinput1 a1[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 a1[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 a1[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 a1[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 a1[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_10_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput6 a1[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_0_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 a1[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 a1[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_0_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19_ net6 _04_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18_ _04_ _05_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor2_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17_ net5 _02_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__and2_1
X_16_ net5 _02_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15_ _03_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14_ _01_ _02_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13_ net2 net1 net3 net4 VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12_ net2 net1 net3 net4 VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11_ net3 _00_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10_ net2 net1 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_5_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

