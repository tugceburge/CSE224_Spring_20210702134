VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO twos_complement
  CLASS BLOCK ;
  FOREIGN twos_complement ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.500 BY 57.120 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 46.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 46.480 ;
    END
  END VPWR
  PIN a1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END a1[0]
  PIN a1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END a1[1]
  PIN a1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END a1[2]
  PIN a1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END a1[3]
  PIN a1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END a1[4]
  PIN a1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END a1[5]
  PIN a1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END a1[6]
  PIN a1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END a1[7]
  PIN b1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END b1[0]
  PIN b1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END b1[1]
  PIN b1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END b1[2]
  PIN b1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END b1[3]
  PIN b1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END b1[4]
  PIN b1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END b1[5]
  PIN b1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END b1[6]
  PIN b1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END b1[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 29.170 46.430 ;
      LAYER li1 ;
        RECT 5.520 10.795 28.980 46.325 ;
      LAYER met1 ;
        RECT 4.210 10.640 28.980 46.480 ;
      LAYER met2 ;
        RECT 4.230 6.955 27.040 48.125 ;
      LAYER met3 ;
        RECT 4.400 47.240 14.610 48.105 ;
        RECT 3.990 45.920 14.610 47.240 ;
        RECT 4.400 44.520 14.610 45.920 ;
        RECT 3.990 43.200 14.610 44.520 ;
        RECT 4.400 41.800 14.610 43.200 ;
        RECT 3.990 40.480 14.610 41.800 ;
        RECT 4.400 39.080 14.610 40.480 ;
        RECT 3.990 37.760 14.610 39.080 ;
        RECT 4.400 36.360 14.610 37.760 ;
        RECT 3.990 35.040 14.610 36.360 ;
        RECT 4.400 33.640 14.610 35.040 ;
        RECT 3.990 32.320 14.610 33.640 ;
        RECT 4.400 30.920 14.610 32.320 ;
        RECT 3.990 29.600 14.610 30.920 ;
        RECT 4.400 28.200 14.610 29.600 ;
        RECT 3.990 26.880 14.610 28.200 ;
        RECT 4.400 25.480 14.610 26.880 ;
        RECT 3.990 24.160 14.610 25.480 ;
        RECT 4.400 22.760 14.610 24.160 ;
        RECT 3.990 21.440 14.610 22.760 ;
        RECT 4.400 20.040 14.610 21.440 ;
        RECT 3.990 18.720 14.610 20.040 ;
        RECT 4.400 17.320 14.610 18.720 ;
        RECT 3.990 16.000 14.610 17.320 ;
        RECT 4.400 14.600 14.610 16.000 ;
        RECT 3.990 13.280 14.610 14.600 ;
        RECT 4.400 11.880 14.610 13.280 ;
        RECT 3.990 10.560 14.610 11.880 ;
        RECT 4.400 9.160 14.610 10.560 ;
        RECT 3.990 7.840 14.610 9.160 ;
        RECT 4.400 6.975 14.610 7.840 ;
  END
END twos_complement
END LIBRARY

