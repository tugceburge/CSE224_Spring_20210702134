magic
tech sky130A
magscale 1 2
timestamp 1745519848
<< nwell >>
rect 1066 2159 5834 9286
<< obsli1 >>
rect 1104 2159 5796 9265
<< obsm1 >>
rect 842 2128 5796 9296
<< obsm2 >>
rect 846 1391 5408 9625
<< metal3 >>
rect 0 9528 800 9648
rect 0 8984 800 9104
rect 0 8440 800 8560
rect 0 7896 800 8016
rect 0 7352 800 7472
rect 0 6808 800 6928
rect 0 6264 800 6384
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 0 4632 800 4752
rect 0 4088 800 4208
rect 0 3544 800 3664
rect 0 3000 800 3120
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 0 1368 800 1488
<< obsm3 >>
rect 880 9448 2922 9621
rect 798 9184 2922 9448
rect 880 8904 2922 9184
rect 798 8640 2922 8904
rect 880 8360 2922 8640
rect 798 8096 2922 8360
rect 880 7816 2922 8096
rect 798 7552 2922 7816
rect 880 7272 2922 7552
rect 798 7008 2922 7272
rect 880 6728 2922 7008
rect 798 6464 2922 6728
rect 880 6184 2922 6464
rect 798 5920 2922 6184
rect 880 5640 2922 5920
rect 798 5376 2922 5640
rect 880 5096 2922 5376
rect 798 4832 2922 5096
rect 880 4552 2922 4832
rect 798 4288 2922 4552
rect 880 4008 2922 4288
rect 798 3744 2922 4008
rect 880 3464 2922 3744
rect 798 3200 2922 3464
rect 880 2920 2922 3200
rect 798 2656 2922 2920
rect 880 2376 2922 2656
rect 798 2112 2922 2376
rect 880 1832 2922 2112
rect 798 1568 2922 1832
rect 880 1395 2922 1568
<< metal4 >>
rect 1944 2128 2264 9296
rect 2604 2128 2924 9296
<< labels >>
rlabel metal4 s 2604 2128 2924 9296 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 9296 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 5176 800 5296 6 a1[0]
port 3 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 a1[1]
port 4 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 a1[2]
port 5 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 a1[3]
port 6 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 a1[4]
port 7 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 a1[5]
port 8 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 a1[6]
port 9 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 a1[7]
port 10 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 b1[0]
port 11 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 b1[1]
port 12 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 b1[2]
port 13 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 b1[3]
port 14 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 b1[4]
port 15 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 b1[5]
port 16 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 b1[6]
port 17 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 b1[7]
port 18 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 6900 11424
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 170272
string GDS_FILE /openlane/designs/twos_complement/runs/RUN_2025.04.24_18.36.13/results/signoff/twos_complement.magic.gds
string GDS_START 83184
<< end >>

